LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.all;
USE  IEEE.STD_LOGIC_ARITH.all;
USE  IEEE.STD_LOGIC_SIGNED.all;


entity LFSR is
	port ( clk, reset : IN std_logic;
		   pipe :	OUT std_logic );
		   
end LSFR;


	